// microprocessor.v

// Generated using ACDS version 15.1 189

`timescale 1 ps / 1 ps
module microprocessor (
		output wire       batharriving_export,    //    batharriving.export
		output wire       bathleaving_export,     //     bathleaving.export
		input  wire       clk_clk,                //             clk.clk
		output wire       drainfinished_export,   //   drainfinished.export
		input  wire       draining_export,        //        draining.export
		output wire       fillfinished_export,    //    fillfinished.export
		input  wire       filling_export,         //         filling.export
		input  wire       innerdoor_export,       //       innerdoor.export
		output wire       innerdoorswitch_export, // innerdoorswitch.export
		input  wire       outerdoor_export,       //       outerdoor.export
		output wire       outerdoorswitch_export, // outerdoorswitch.export
		output wire       personcheck_export,     //     personcheck.export
		output wire       pressurecheck_export,   //   pressurecheck.export
		input  wire       reset_reset_n,          //           reset.reset_n
		input  wire [3:0] resetleds_export,       //       resetleds.export
		output wire       waitfinished_export,    //    waitfinished.export
		input  wire       waiting_export          //         waiting.export
	);

	wire  [31:0] nios2_processor_data_master_readdata;                          // mm_interconnect_0:nios2_processor_data_master_readdata -> nios2_processor:d_readdata
	wire         nios2_processor_data_master_waitrequest;                       // mm_interconnect_0:nios2_processor_data_master_waitrequest -> nios2_processor:d_waitrequest
	wire         nios2_processor_data_master_debugaccess;                       // nios2_processor:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_processor_data_master_debugaccess
	wire  [13:0] nios2_processor_data_master_address;                           // nios2_processor:d_address -> mm_interconnect_0:nios2_processor_data_master_address
	wire   [3:0] nios2_processor_data_master_byteenable;                        // nios2_processor:d_byteenable -> mm_interconnect_0:nios2_processor_data_master_byteenable
	wire         nios2_processor_data_master_read;                              // nios2_processor:d_read -> mm_interconnect_0:nios2_processor_data_master_read
	wire         nios2_processor_data_master_write;                             // nios2_processor:d_write -> mm_interconnect_0:nios2_processor_data_master_write
	wire  [31:0] nios2_processor_data_master_writedata;                         // nios2_processor:d_writedata -> mm_interconnect_0:nios2_processor_data_master_writedata
	wire  [31:0] nios2_processor_instruction_master_readdata;                   // mm_interconnect_0:nios2_processor_instruction_master_readdata -> nios2_processor:i_readdata
	wire         nios2_processor_instruction_master_waitrequest;                // mm_interconnect_0:nios2_processor_instruction_master_waitrequest -> nios2_processor:i_waitrequest
	wire  [13:0] nios2_processor_instruction_master_address;                    // nios2_processor:i_address -> mm_interconnect_0:nios2_processor_instruction_master_address
	wire         nios2_processor_instruction_master_read;                       // nios2_processor:i_read -> mm_interconnect_0:nios2_processor_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;        // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;     // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_processor_debug_mem_slave_readdata;    // nios2_processor:debug_mem_slave_readdata -> mm_interconnect_0:nios2_processor_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_waitrequest; // nios2_processor:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_processor_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_processor_debug_mem_slave_debugaccess -> nios2_processor:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_processor_debug_mem_slave_address;     // mm_interconnect_0:nios2_processor_debug_mem_slave_address -> nios2_processor:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_read;        // mm_interconnect_0:nios2_processor_debug_mem_slave_read -> nios2_processor:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_processor_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_processor_debug_mem_slave_byteenable -> nios2_processor:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_write;       // mm_interconnect_0:nios2_processor_debug_mem_slave_write -> nios2_processor:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_processor_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_processor_debug_mem_slave_writedata -> nios2_processor:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                 // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                   // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory_s1_address;                    // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                 // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                      // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                  // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                      // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire  [31:0] mm_interconnect_0_filling_s1_readdata;                         // Filling:readdata -> mm_interconnect_0:Filling_s1_readdata
	wire   [1:0] mm_interconnect_0_filling_s1_address;                          // mm_interconnect_0:Filling_s1_address -> Filling:address
	wire  [31:0] mm_interconnect_0_draining_s1_readdata;                        // Draining:readdata -> mm_interconnect_0:Draining_s1_readdata
	wire   [1:0] mm_interconnect_0_draining_s1_address;                         // mm_interconnect_0:Draining_s1_address -> Draining:address
	wire  [31:0] mm_interconnect_0_innerdoor_s1_readdata;                       // innerDoor:readdata -> mm_interconnect_0:innerDoor_s1_readdata
	wire   [1:0] mm_interconnect_0_innerdoor_s1_address;                        // mm_interconnect_0:innerDoor_s1_address -> innerDoor:address
	wire  [31:0] mm_interconnect_0_outerdoor_s1_readdata;                       // outerDoor:readdata -> mm_interconnect_0:outerDoor_s1_readdata
	wire   [1:0] mm_interconnect_0_outerdoor_s1_address;                        // mm_interconnect_0:outerDoor_s1_address -> outerDoor:address
	wire  [31:0] mm_interconnect_0_resetleds_s1_readdata;                       // resetLeds:readdata -> mm_interconnect_0:resetLeds_s1_readdata
	wire   [1:0] mm_interconnect_0_resetleds_s1_address;                        // mm_interconnect_0:resetLeds_s1_address -> resetLeds:address
	wire         mm_interconnect_0_bathleaving_s1_chipselect;                   // mm_interconnect_0:bathLeaving_s1_chipselect -> bathLeaving:chipselect
	wire  [31:0] mm_interconnect_0_bathleaving_s1_readdata;                     // bathLeaving:readdata -> mm_interconnect_0:bathLeaving_s1_readdata
	wire   [1:0] mm_interconnect_0_bathleaving_s1_address;                      // mm_interconnect_0:bathLeaving_s1_address -> bathLeaving:address
	wire         mm_interconnect_0_bathleaving_s1_write;                        // mm_interconnect_0:bathLeaving_s1_write -> bathLeaving:write_n
	wire  [31:0] mm_interconnect_0_bathleaving_s1_writedata;                    // mm_interconnect_0:bathLeaving_s1_writedata -> bathLeaving:writedata
	wire         mm_interconnect_0_batharriving_s1_chipselect;                  // mm_interconnect_0:bathArriving_s1_chipselect -> bathArriving:chipselect
	wire  [31:0] mm_interconnect_0_batharriving_s1_readdata;                    // bathArriving:readdata -> mm_interconnect_0:bathArriving_s1_readdata
	wire   [1:0] mm_interconnect_0_batharriving_s1_address;                     // mm_interconnect_0:bathArriving_s1_address -> bathArriving:address
	wire         mm_interconnect_0_batharriving_s1_write;                       // mm_interconnect_0:bathArriving_s1_write -> bathArriving:write_n
	wire  [31:0] mm_interconnect_0_batharriving_s1_writedata;                   // mm_interconnect_0:bathArriving_s1_writedata -> bathArriving:writedata
	wire         mm_interconnect_0_personcheck_s1_chipselect;                   // mm_interconnect_0:personCheck_s1_chipselect -> personCheck:chipselect
	wire  [31:0] mm_interconnect_0_personcheck_s1_readdata;                     // personCheck:readdata -> mm_interconnect_0:personCheck_s1_readdata
	wire   [1:0] mm_interconnect_0_personcheck_s1_address;                      // mm_interconnect_0:personCheck_s1_address -> personCheck:address
	wire         mm_interconnect_0_personcheck_s1_write;                        // mm_interconnect_0:personCheck_s1_write -> personCheck:write_n
	wire  [31:0] mm_interconnect_0_personcheck_s1_writedata;                    // mm_interconnect_0:personCheck_s1_writedata -> personCheck:writedata
	wire         mm_interconnect_0_pressurecheck_s1_chipselect;                 // mm_interconnect_0:pressureCheck_s1_chipselect -> pressureCheck:chipselect
	wire  [31:0] mm_interconnect_0_pressurecheck_s1_readdata;                   // pressureCheck:readdata -> mm_interconnect_0:pressureCheck_s1_readdata
	wire   [1:0] mm_interconnect_0_pressurecheck_s1_address;                    // mm_interconnect_0:pressureCheck_s1_address -> pressureCheck:address
	wire         mm_interconnect_0_pressurecheck_s1_write;                      // mm_interconnect_0:pressureCheck_s1_write -> pressureCheck:write_n
	wire  [31:0] mm_interconnect_0_pressurecheck_s1_writedata;                  // mm_interconnect_0:pressureCheck_s1_writedata -> pressureCheck:writedata
	wire         mm_interconnect_0_innerdoorswitch_s1_chipselect;               // mm_interconnect_0:innerDoorSwitch_s1_chipselect -> innerDoorSwitch:chipselect
	wire  [31:0] mm_interconnect_0_innerdoorswitch_s1_readdata;                 // innerDoorSwitch:readdata -> mm_interconnect_0:innerDoorSwitch_s1_readdata
	wire   [1:0] mm_interconnect_0_innerdoorswitch_s1_address;                  // mm_interconnect_0:innerDoorSwitch_s1_address -> innerDoorSwitch:address
	wire         mm_interconnect_0_innerdoorswitch_s1_write;                    // mm_interconnect_0:innerDoorSwitch_s1_write -> innerDoorSwitch:write_n
	wire  [31:0] mm_interconnect_0_innerdoorswitch_s1_writedata;                // mm_interconnect_0:innerDoorSwitch_s1_writedata -> innerDoorSwitch:writedata
	wire         mm_interconnect_0_outerdoorswitch_s1_chipselect;               // mm_interconnect_0:outerDoorSwitch_s1_chipselect -> outerDoorSwitch:chipselect
	wire  [31:0] mm_interconnect_0_outerdoorswitch_s1_readdata;                 // outerDoorSwitch:readdata -> mm_interconnect_0:outerDoorSwitch_s1_readdata
	wire   [1:0] mm_interconnect_0_outerdoorswitch_s1_address;                  // mm_interconnect_0:outerDoorSwitch_s1_address -> outerDoorSwitch:address
	wire         mm_interconnect_0_outerdoorswitch_s1_write;                    // mm_interconnect_0:outerDoorSwitch_s1_write -> outerDoorSwitch:write_n
	wire  [31:0] mm_interconnect_0_outerdoorswitch_s1_writedata;                // mm_interconnect_0:outerDoorSwitch_s1_writedata -> outerDoorSwitch:writedata
	wire         mm_interconnect_0_drainfinished_s1_chipselect;                 // mm_interconnect_0:drainFinished_s1_chipselect -> drainFinished:chipselect
	wire  [31:0] mm_interconnect_0_drainfinished_s1_readdata;                   // drainFinished:readdata -> mm_interconnect_0:drainFinished_s1_readdata
	wire   [1:0] mm_interconnect_0_drainfinished_s1_address;                    // mm_interconnect_0:drainFinished_s1_address -> drainFinished:address
	wire         mm_interconnect_0_drainfinished_s1_write;                      // mm_interconnect_0:drainFinished_s1_write -> drainFinished:write_n
	wire  [31:0] mm_interconnect_0_drainfinished_s1_writedata;                  // mm_interconnect_0:drainFinished_s1_writedata -> drainFinished:writedata
	wire         mm_interconnect_0_fillfinished_s1_chipselect;                  // mm_interconnect_0:fillFinished_s1_chipselect -> fillFinished:chipselect
	wire  [31:0] mm_interconnect_0_fillfinished_s1_readdata;                    // fillFinished:readdata -> mm_interconnect_0:fillFinished_s1_readdata
	wire   [1:0] mm_interconnect_0_fillfinished_s1_address;                     // mm_interconnect_0:fillFinished_s1_address -> fillFinished:address
	wire         mm_interconnect_0_fillfinished_s1_write;                       // mm_interconnect_0:fillFinished_s1_write -> fillFinished:write_n
	wire  [31:0] mm_interconnect_0_fillfinished_s1_writedata;                   // mm_interconnect_0:fillFinished_s1_writedata -> fillFinished:writedata
	wire         mm_interconnect_0_waitfinished_s1_chipselect;                  // mm_interconnect_0:waitFinished_s1_chipselect -> waitFinished:chipselect
	wire  [31:0] mm_interconnect_0_waitfinished_s1_readdata;                    // waitFinished:readdata -> mm_interconnect_0:waitFinished_s1_readdata
	wire   [1:0] mm_interconnect_0_waitfinished_s1_address;                     // mm_interconnect_0:waitFinished_s1_address -> waitFinished:address
	wire         mm_interconnect_0_waitfinished_s1_write;                       // mm_interconnect_0:waitFinished_s1_write -> waitFinished:write_n
	wire  [31:0] mm_interconnect_0_waitfinished_s1_writedata;                   // mm_interconnect_0:waitFinished_s1_writedata -> waitFinished:writedata
	wire  [31:0] mm_interconnect_0_waiting_s1_readdata;                         // waiting:readdata -> mm_interconnect_0:waiting_s1_readdata
	wire   [1:0] mm_interconnect_0_waiting_s1_address;                          // mm_interconnect_0:waiting_s1_address -> waiting:address
	wire         irq_mapper_receiver0_irq;                                      // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_processor_irq_irq;                                       // irq_mapper:sender_irq -> nios2_processor:irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [Draining:reset_n, Filling:reset_n, bathArriving:reset_n, bathLeaving:reset_n, drainFinished:reset_n, fillFinished:reset_n, innerDoor:reset_n, innerDoorSwitch:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_processor_reset_reset_bridge_in_reset_reset, nios2_processor:reset_n, onchip_memory:reset, outerDoor:reset_n, outerDoorSwitch:reset_n, personCheck:reset_n, pressureCheck:reset_n, resetLeds:reset_n, rst_translator:in_reset, waitFinished:reset_n, waiting:reset_n]
	wire         rst_controller_reset_out_reset_req;                            // rst_controller:reset_req -> [nios2_processor:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios2_processor_debug_reset_request_reset;                     // nios2_processor:debug_reset_request -> rst_controller:reset_in1

	microprocessor_Draining draining (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_draining_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_draining_s1_readdata), //                    .readdata
		.in_port  (draining_export)                         // external_connection.export
	);

	microprocessor_Draining filling (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_filling_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_filling_s1_readdata), //                    .readdata
		.in_port  (filling_export)                         // external_connection.export
	);

	microprocessor_bathArriving batharriving (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_batharriving_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_batharriving_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_batharriving_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_batharriving_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_batharriving_s1_readdata),   //                    .readdata
		.out_port   (batharriving_export)                           // external_connection.export
	);

	microprocessor_bathArriving bathleaving (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_bathleaving_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bathleaving_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bathleaving_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bathleaving_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bathleaving_s1_readdata),   //                    .readdata
		.out_port   (bathleaving_export)                           // external_connection.export
	);

	microprocessor_bathArriving drainfinished (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_drainfinished_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_drainfinished_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_drainfinished_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_drainfinished_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_drainfinished_s1_readdata),   //                    .readdata
		.out_port   (drainfinished_export)                           // external_connection.export
	);

	microprocessor_bathArriving fillfinished (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_fillfinished_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fillfinished_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fillfinished_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fillfinished_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fillfinished_s1_readdata),   //                    .readdata
		.out_port   (fillfinished_export)                           // external_connection.export
	);

	microprocessor_Draining innerdoor (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_innerdoor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_innerdoor_s1_readdata), //                    .readdata
		.in_port  (innerdoor_export)                         // external_connection.export
	);

	microprocessor_bathArriving innerdoorswitch (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_innerdoorswitch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_innerdoorswitch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_innerdoorswitch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_innerdoorswitch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_innerdoorswitch_s1_readdata),   //                    .readdata
		.out_port   (innerdoorswitch_export)                           // external_connection.export
	);

	microprocessor_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	microprocessor_nios2_processor nios2_processor (
		.clk                                 (clk_clk),                                                       //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                               //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                            //                          .reset_req
		.d_address                           (nios2_processor_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_processor_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_processor_data_master_read),                              //                          .read
		.d_readdata                          (nios2_processor_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_processor_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_processor_data_master_write),                             //                          .write
		.d_writedata                         (nios2_processor_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_processor_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_processor_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_processor_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_processor_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_processor_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_processor_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_processor_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_processor_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_processor_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_processor_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_processor_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_processor_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_processor_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_processor_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                               // custom_instruction_master.readra
	);

	microprocessor_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	microprocessor_Draining outerdoor (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_outerdoor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_outerdoor_s1_readdata), //                    .readdata
		.in_port  (outerdoor_export)                         // external_connection.export
	);

	microprocessor_bathArriving outerdoorswitch (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_outerdoorswitch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_outerdoorswitch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_outerdoorswitch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_outerdoorswitch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_outerdoorswitch_s1_readdata),   //                    .readdata
		.out_port   (outerdoorswitch_export)                           // external_connection.export
	);

	microprocessor_bathArriving personcheck (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_personcheck_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_personcheck_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_personcheck_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_personcheck_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_personcheck_s1_readdata),   //                    .readdata
		.out_port   (personcheck_export)                           // external_connection.export
	);

	microprocessor_bathArriving pressurecheck (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pressurecheck_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pressurecheck_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pressurecheck_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pressurecheck_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pressurecheck_s1_readdata),   //                    .readdata
		.out_port   (pressurecheck_export)                           // external_connection.export
	);

	microprocessor_resetLeds resetleds (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_resetleds_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_resetleds_s1_readdata), //                    .readdata
		.in_port  (resetleds_export)                         // external_connection.export
	);

	microprocessor_bathArriving waitfinished (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_waitfinished_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_waitfinished_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_waitfinished_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_waitfinished_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_waitfinished_s1_readdata),   //                    .readdata
		.out_port   (waitfinished_export)                           // external_connection.export
	);

	microprocessor_Draining waiting (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_waiting_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_waiting_s1_readdata), //                    .readdata
		.in_port  (waiting_export)                         // external_connection.export
	);

	microprocessor_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                     (clk_clk),                                                       //                                   clk_0_clk.clk
		.nios2_processor_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // nios2_processor_reset_reset_bridge_in_reset.reset
		.nios2_processor_data_master_address               (nios2_processor_data_master_address),                           //                 nios2_processor_data_master.address
		.nios2_processor_data_master_waitrequest           (nios2_processor_data_master_waitrequest),                       //                                            .waitrequest
		.nios2_processor_data_master_byteenable            (nios2_processor_data_master_byteenable),                        //                                            .byteenable
		.nios2_processor_data_master_read                  (nios2_processor_data_master_read),                              //                                            .read
		.nios2_processor_data_master_readdata              (nios2_processor_data_master_readdata),                          //                                            .readdata
		.nios2_processor_data_master_write                 (nios2_processor_data_master_write),                             //                                            .write
		.nios2_processor_data_master_writedata             (nios2_processor_data_master_writedata),                         //                                            .writedata
		.nios2_processor_data_master_debugaccess           (nios2_processor_data_master_debugaccess),                       //                                            .debugaccess
		.nios2_processor_instruction_master_address        (nios2_processor_instruction_master_address),                    //          nios2_processor_instruction_master.address
		.nios2_processor_instruction_master_waitrequest    (nios2_processor_instruction_master_waitrequest),                //                                            .waitrequest
		.nios2_processor_instruction_master_read           (nios2_processor_instruction_master_read),                       //                                            .read
		.nios2_processor_instruction_master_readdata       (nios2_processor_instruction_master_readdata),                   //                                            .readdata
		.bathArriving_s1_address                           (mm_interconnect_0_batharriving_s1_address),                     //                             bathArriving_s1.address
		.bathArriving_s1_write                             (mm_interconnect_0_batharriving_s1_write),                       //                                            .write
		.bathArriving_s1_readdata                          (mm_interconnect_0_batharriving_s1_readdata),                    //                                            .readdata
		.bathArriving_s1_writedata                         (mm_interconnect_0_batharriving_s1_writedata),                   //                                            .writedata
		.bathArriving_s1_chipselect                        (mm_interconnect_0_batharriving_s1_chipselect),                  //                                            .chipselect
		.bathLeaving_s1_address                            (mm_interconnect_0_bathleaving_s1_address),                      //                              bathLeaving_s1.address
		.bathLeaving_s1_write                              (mm_interconnect_0_bathleaving_s1_write),                        //                                            .write
		.bathLeaving_s1_readdata                           (mm_interconnect_0_bathleaving_s1_readdata),                     //                                            .readdata
		.bathLeaving_s1_writedata                          (mm_interconnect_0_bathleaving_s1_writedata),                    //                                            .writedata
		.bathLeaving_s1_chipselect                         (mm_interconnect_0_bathleaving_s1_chipselect),                   //                                            .chipselect
		.drainFinished_s1_address                          (mm_interconnect_0_drainfinished_s1_address),                    //                            drainFinished_s1.address
		.drainFinished_s1_write                            (mm_interconnect_0_drainfinished_s1_write),                      //                                            .write
		.drainFinished_s1_readdata                         (mm_interconnect_0_drainfinished_s1_readdata),                   //                                            .readdata
		.drainFinished_s1_writedata                        (mm_interconnect_0_drainfinished_s1_writedata),                  //                                            .writedata
		.drainFinished_s1_chipselect                       (mm_interconnect_0_drainfinished_s1_chipselect),                 //                                            .chipselect
		.Draining_s1_address                               (mm_interconnect_0_draining_s1_address),                         //                                 Draining_s1.address
		.Draining_s1_readdata                              (mm_interconnect_0_draining_s1_readdata),                        //                                            .readdata
		.fillFinished_s1_address                           (mm_interconnect_0_fillfinished_s1_address),                     //                             fillFinished_s1.address
		.fillFinished_s1_write                             (mm_interconnect_0_fillfinished_s1_write),                       //                                            .write
		.fillFinished_s1_readdata                          (mm_interconnect_0_fillfinished_s1_readdata),                    //                                            .readdata
		.fillFinished_s1_writedata                         (mm_interconnect_0_fillfinished_s1_writedata),                   //                                            .writedata
		.fillFinished_s1_chipselect                        (mm_interconnect_0_fillfinished_s1_chipselect),                  //                                            .chipselect
		.Filling_s1_address                                (mm_interconnect_0_filling_s1_address),                          //                                  Filling_s1.address
		.Filling_s1_readdata                               (mm_interconnect_0_filling_s1_readdata),                         //                                            .readdata
		.innerDoor_s1_address                              (mm_interconnect_0_innerdoor_s1_address),                        //                                innerDoor_s1.address
		.innerDoor_s1_readdata                             (mm_interconnect_0_innerdoor_s1_readdata),                       //                                            .readdata
		.innerDoorSwitch_s1_address                        (mm_interconnect_0_innerdoorswitch_s1_address),                  //                          innerDoorSwitch_s1.address
		.innerDoorSwitch_s1_write                          (mm_interconnect_0_innerdoorswitch_s1_write),                    //                                            .write
		.innerDoorSwitch_s1_readdata                       (mm_interconnect_0_innerdoorswitch_s1_readdata),                 //                                            .readdata
		.innerDoorSwitch_s1_writedata                      (mm_interconnect_0_innerdoorswitch_s1_writedata),                //                                            .writedata
		.innerDoorSwitch_s1_chipselect                     (mm_interconnect_0_innerdoorswitch_s1_chipselect),               //                                            .chipselect
		.jtag_uart_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),         //                 jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),           //                                            .write
		.jtag_uart_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),            //                                            .read
		.jtag_uart_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),        //                                            .readdata
		.jtag_uart_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),       //                                            .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),     //                                            .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),      //                                            .chipselect
		.nios2_processor_debug_mem_slave_address           (mm_interconnect_0_nios2_processor_debug_mem_slave_address),     //             nios2_processor_debug_mem_slave.address
		.nios2_processor_debug_mem_slave_write             (mm_interconnect_0_nios2_processor_debug_mem_slave_write),       //                                            .write
		.nios2_processor_debug_mem_slave_read              (mm_interconnect_0_nios2_processor_debug_mem_slave_read),        //                                            .read
		.nios2_processor_debug_mem_slave_readdata          (mm_interconnect_0_nios2_processor_debug_mem_slave_readdata),    //                                            .readdata
		.nios2_processor_debug_mem_slave_writedata         (mm_interconnect_0_nios2_processor_debug_mem_slave_writedata),   //                                            .writedata
		.nios2_processor_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_processor_debug_mem_slave_byteenable),  //                                            .byteenable
		.nios2_processor_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_processor_debug_mem_slave_waitrequest), //                                            .waitrequest
		.nios2_processor_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_processor_debug_mem_slave_debugaccess), //                                            .debugaccess
		.onchip_memory_s1_address                          (mm_interconnect_0_onchip_memory_s1_address),                    //                            onchip_memory_s1.address
		.onchip_memory_s1_write                            (mm_interconnect_0_onchip_memory_s1_write),                      //                                            .write
		.onchip_memory_s1_readdata                         (mm_interconnect_0_onchip_memory_s1_readdata),                   //                                            .readdata
		.onchip_memory_s1_writedata                        (mm_interconnect_0_onchip_memory_s1_writedata),                  //                                            .writedata
		.onchip_memory_s1_byteenable                       (mm_interconnect_0_onchip_memory_s1_byteenable),                 //                                            .byteenable
		.onchip_memory_s1_chipselect                       (mm_interconnect_0_onchip_memory_s1_chipselect),                 //                                            .chipselect
		.onchip_memory_s1_clken                            (mm_interconnect_0_onchip_memory_s1_clken),                      //                                            .clken
		.outerDoor_s1_address                              (mm_interconnect_0_outerdoor_s1_address),                        //                                outerDoor_s1.address
		.outerDoor_s1_readdata                             (mm_interconnect_0_outerdoor_s1_readdata),                       //                                            .readdata
		.outerDoorSwitch_s1_address                        (mm_interconnect_0_outerdoorswitch_s1_address),                  //                          outerDoorSwitch_s1.address
		.outerDoorSwitch_s1_write                          (mm_interconnect_0_outerdoorswitch_s1_write),                    //                                            .write
		.outerDoorSwitch_s1_readdata                       (mm_interconnect_0_outerdoorswitch_s1_readdata),                 //                                            .readdata
		.outerDoorSwitch_s1_writedata                      (mm_interconnect_0_outerdoorswitch_s1_writedata),                //                                            .writedata
		.outerDoorSwitch_s1_chipselect                     (mm_interconnect_0_outerdoorswitch_s1_chipselect),               //                                            .chipselect
		.personCheck_s1_address                            (mm_interconnect_0_personcheck_s1_address),                      //                              personCheck_s1.address
		.personCheck_s1_write                              (mm_interconnect_0_personcheck_s1_write),                        //                                            .write
		.personCheck_s1_readdata                           (mm_interconnect_0_personcheck_s1_readdata),                     //                                            .readdata
		.personCheck_s1_writedata                          (mm_interconnect_0_personcheck_s1_writedata),                    //                                            .writedata
		.personCheck_s1_chipselect                         (mm_interconnect_0_personcheck_s1_chipselect),                   //                                            .chipselect
		.pressureCheck_s1_address                          (mm_interconnect_0_pressurecheck_s1_address),                    //                            pressureCheck_s1.address
		.pressureCheck_s1_write                            (mm_interconnect_0_pressurecheck_s1_write),                      //                                            .write
		.pressureCheck_s1_readdata                         (mm_interconnect_0_pressurecheck_s1_readdata),                   //                                            .readdata
		.pressureCheck_s1_writedata                        (mm_interconnect_0_pressurecheck_s1_writedata),                  //                                            .writedata
		.pressureCheck_s1_chipselect                       (mm_interconnect_0_pressurecheck_s1_chipselect),                 //                                            .chipselect
		.resetLeds_s1_address                              (mm_interconnect_0_resetleds_s1_address),                        //                                resetLeds_s1.address
		.resetLeds_s1_readdata                             (mm_interconnect_0_resetleds_s1_readdata),                       //                                            .readdata
		.waitFinished_s1_address                           (mm_interconnect_0_waitfinished_s1_address),                     //                             waitFinished_s1.address
		.waitFinished_s1_write                             (mm_interconnect_0_waitfinished_s1_write),                       //                                            .write
		.waitFinished_s1_readdata                          (mm_interconnect_0_waitfinished_s1_readdata),                    //                                            .readdata
		.waitFinished_s1_writedata                         (mm_interconnect_0_waitfinished_s1_writedata),                   //                                            .writedata
		.waitFinished_s1_chipselect                        (mm_interconnect_0_waitfinished_s1_chipselect),                  //                                            .chipselect
		.waiting_s1_address                                (mm_interconnect_0_waiting_s1_address),                          //                                  waiting_s1.address
		.waiting_s1_readdata                               (mm_interconnect_0_waiting_s1_readdata)                          //                                            .readdata
	);

	microprocessor_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_processor_irq_irq)         //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                            // reset_in0.reset
		.reset_in1      (nios2_processor_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                   //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),            // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),        //          .reset_req
		.reset_req_in0  (1'b0),                                      // (terminated)
		.reset_req_in1  (1'b0),                                      // (terminated)
		.reset_in2      (1'b0),                                      // (terminated)
		.reset_req_in2  (1'b0),                                      // (terminated)
		.reset_in3      (1'b0),                                      // (terminated)
		.reset_req_in3  (1'b0),                                      // (terminated)
		.reset_in4      (1'b0),                                      // (terminated)
		.reset_req_in4  (1'b0),                                      // (terminated)
		.reset_in5      (1'b0),                                      // (terminated)
		.reset_req_in5  (1'b0),                                      // (terminated)
		.reset_in6      (1'b0),                                      // (terminated)
		.reset_req_in6  (1'b0),                                      // (terminated)
		.reset_in7      (1'b0),                                      // (terminated)
		.reset_req_in7  (1'b0),                                      // (terminated)
		.reset_in8      (1'b0),                                      // (terminated)
		.reset_req_in8  (1'b0),                                      // (terminated)
		.reset_in9      (1'b0),                                      // (terminated)
		.reset_req_in9  (1'b0),                                      // (terminated)
		.reset_in10     (1'b0),                                      // (terminated)
		.reset_req_in10 (1'b0),                                      // (terminated)
		.reset_in11     (1'b0),                                      // (terminated)
		.reset_req_in11 (1'b0),                                      // (terminated)
		.reset_in12     (1'b0),                                      // (terminated)
		.reset_req_in12 (1'b0),                                      // (terminated)
		.reset_in13     (1'b0),                                      // (terminated)
		.reset_req_in13 (1'b0),                                      // (terminated)
		.reset_in14     (1'b0),                                      // (terminated)
		.reset_req_in14 (1'b0),                                      // (terminated)
		.reset_in15     (1'b0),                                      // (terminated)
		.reset_req_in15 (1'b0)                                       // (terminated)
	);

endmodule
